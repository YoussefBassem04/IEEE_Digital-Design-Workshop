module and_gate (input A,B,output out);

assign out = A && B;



endmodule