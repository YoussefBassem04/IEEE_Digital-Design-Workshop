module Half_Adder(input A,B, output s,c);

assign {c,s} = A + B;


endmodule